--F Function of SHA-3
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;	
