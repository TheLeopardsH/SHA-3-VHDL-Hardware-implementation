library ieee;
use ieee.std_logic_1164.all;

package keccakVar is

	constant i : integer :=5;
	constant j : integer :=5;
	constant k : integer :=64;
	
	type array1D is array((k-1) downto 0) of std_logic;
	type array2D is array((j-1) downto 0) of array1D ;
	type array3D_state is array((i-1) downto 0) of array2D ;
	
end package;
